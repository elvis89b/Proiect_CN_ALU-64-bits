library verilog;
use verilog.vl_types.all;
entity ml_csea_8_tb is
end ml_csea_8_tb;
