library verilog;
use verilog.vl_types.all;
entity bitwise_xnor_tb is
end bitwise_xnor_tb;
