library verilog;
use verilog.vl_types.all;
entity mux8to1_tb is
end mux8to1_tb;
