library verilog;
use verilog.vl_types.all;
entity sh_reg_tb is
end sh_reg_tb;
