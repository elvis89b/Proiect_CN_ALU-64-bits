library verilog;
use verilog.vl_types.all;
entity bitwise_nor_tb is
end bitwise_nor_tb;
