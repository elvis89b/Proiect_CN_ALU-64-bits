library verilog;
use verilog.vl_types.all;
entity rotl_tb is
end rotl_tb;
