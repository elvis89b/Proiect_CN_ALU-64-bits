library verilog;
use verilog.vl_types.all;
entity srl_tb is
end srl_tb;
