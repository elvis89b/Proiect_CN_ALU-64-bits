module bitwise_or (
  input in_0,
  input in_1,
  output or_
);

  assign or_ = in_0 | in_1;
  
endmodule