library verilog;
use verilog.vl_types.all;
entity substractor_tb is
end substractor_tb;
