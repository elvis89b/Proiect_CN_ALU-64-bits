library verilog;
use verilog.vl_types.all;
entity mux2to1_tb is
end mux2to1_tb;
