library verilog;
use verilog.vl_types.all;
entity not_wordgate_tb is
end not_wordgate_tb;
