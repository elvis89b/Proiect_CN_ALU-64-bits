library verilog;
use verilog.vl_types.all;
entity bitwise_not_tb is
end bitwise_not_tb;
