library verilog;
use verilog.vl_types.all;
entity shift_rotate_unit_tb is
end shift_rotate_unit_tb;
