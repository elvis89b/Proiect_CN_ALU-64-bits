library verilog;
use verilog.vl_types.all;
entity xor_wordgate_tb is
end xor_wordgate_tb;
