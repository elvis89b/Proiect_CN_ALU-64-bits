library verilog;
use verilog.vl_types.all;
entity or_wordgate_tb is
end or_wordgate_tb;
