library verilog;
use verilog.vl_types.all;
entity sll_tb is
end sll_tb;
