module bitwise_xor (
  input in_0,
  input in_1,
  output xor_
);

  assign xor_ = in_0 ^ in_1;
  
endmodule