library verilog;
use verilog.vl_types.all;
entity ALU_64_tb is
end ALU_64_tb;
