library verilog;
use verilog.vl_types.all;
entity br2_tb is
end br2_tb;
