library verilog;
use verilog.vl_types.all;
entity sra_tb is
end sra_tb;
