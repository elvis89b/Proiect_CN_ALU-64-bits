library verilog;
use verilog.vl_types.all;
entity reg_M_tb is
end reg_M_tb;
