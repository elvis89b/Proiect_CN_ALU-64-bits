library verilog;
use verilog.vl_types.all;
entity nand_wordgate_tb is
end nand_wordgate_tb;
