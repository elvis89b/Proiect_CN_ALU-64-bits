library verilog;
use verilog.vl_types.all;
entity reg_A_tb is
end reg_A_tb;
