library verilog;
use verilog.vl_types.all;
entity bitwise_xor_tb is
end bitwise_xor_tb;
