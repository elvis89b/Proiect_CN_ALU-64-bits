library verilog;
use verilog.vl_types.all;
entity bitwise_nand_tb is
end bitwise_nand_tb;
