module bitwise_not (
  input in,
  output not_
);

  assign not_ = ~in;
  
endmodule