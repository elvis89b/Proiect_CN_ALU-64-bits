library verilog;
use verilog.vl_types.all;
entity mux16to1_tb is
end mux16to1_tb;
