library verilog;
use verilog.vl_types.all;
entity xnor_wordgate_tb is
end xnor_wordgate_tb;
