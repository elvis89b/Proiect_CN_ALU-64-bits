library verilog;
use verilog.vl_types.all;
entity reg_Q_tb is
end reg_Q_tb;
