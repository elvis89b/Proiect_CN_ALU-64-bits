library verilog;
use verilog.vl_types.all;
entity bitwise_or_tb is
end bitwise_or_tb;
