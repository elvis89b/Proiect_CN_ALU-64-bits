library verilog;
use verilog.vl_types.all;
entity csea_level_tb is
end csea_level_tb;
