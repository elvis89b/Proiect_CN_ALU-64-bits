library verilog;
use verilog.vl_types.all;
entity logic_unit_tb is
end logic_unit_tb;
