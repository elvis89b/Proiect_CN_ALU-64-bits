library verilog;
use verilog.vl_types.all;
entity rotr_tb is
end rotr_tb;
