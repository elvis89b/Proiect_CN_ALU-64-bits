library verilog;
use verilog.vl_types.all;
entity nor_wordgate_tb is
end nor_wordgate_tb;
