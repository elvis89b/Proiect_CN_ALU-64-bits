library verilog;
use verilog.vl_types.all;
entity sla_tb is
end sla_tb;
